library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;
use ieee.math_real.all;

entity Instruction_Memory is
  port(  read_ena : in std_logic;
         address : in std_logic_vector(15 downto 0);
			instruction_out  : out std_logic_vector(15 downto 0):= (others=> 'X'));
end Instruction_Memory;

architecture Instruction_behave of Instruction_Memory is
type memory_table is array ( 255 downto 0) of std_logic_vector(15 downto 0);
signal i_memory: memory_table :=(

                                 

											0 =>"0011000000000000",----------------------------LHI -Load R0 with 0
                                 1 =>"0011001000000001",----------------------------LHI -Load R1 with 128
											2 =>"0011010000000010",----------------------------LHI -Load R2 with 256
											3 =>"0011011000000011",----------------------------LHI -Load R3 with 384
											4 =>"0011100000000100",----------------------------LHI -Load R4 with 512
											5 =>"0011101000000101",----------------------------LHI -Load R5 with 640
											6 =>"0011110000000110",----------------------------LHI -Load R6 with 768
											
											7 =>"0001001001010000",----------------------------ADD(r2=r1 + r1)
											8 =>"0011111000000111",----------------------------LHI -Load R7 with 896
											9 =>"0011111000000111",----------------------------LHI -Load R7 with 896
											10=>"0101001001000000",----------------------------SW - Load memory address(128) with 128
											11=>"0011110000000110",----------------------------LHI -Load R6 with 768
											12 =>"0001000001010010",----------------------------ADC(r2=r1+r0)
                                 13 =>"0011111000000111",----------------------------LHI -Load R7 with 896
											14 => "0100000001000000",----------------------------LW  -Load R1 with 128
											
								
     										15=>"0001001010010000",----------------------------r2=r1+r2
											
--											9 =>"0001000001010000",----------------------------ADD -Load R2 with 128(R2=R0+R1)
										 
										 
--											10=>"0101001001000000",----------------------------SW - Load memory address(128) with 128
--											11=>"0101010000000000",----------------------------SW - Load memory address(0) with 256 
--											12=>"0011111000000101",----------------------------LHI -Load R7 with 640
--											13=>"0011111000000001",----------------------------LHI -Load R7 with 128
--											14=>"0100010010000000",----------------------------LW  -Load R2 with 256
--											15=>"0001000001010010",----------------------------ADC -do not Load R2 with 16(because carry_flag is 0)
--											16=>"0001000001010001",----------------------------ADZ -do not Load R2 with 16(because zero_flag is 0)
--											17=>"0001000001010011",----------------------------ADL -Load R2 with 32
--											18=>"0010000001010000",----------------------------NDU 
--											19=>"0010000001010010",----------------------------NDC 
--											20=>"0010000001010001",----------------------------NDZ 
--											21=>"0011010000000010",----------------------------LHI -Load R2 with 256
--											22=>"1000110111001000",--beq to 30
--											23=>"0011011000000010",----------------------------LHI -Load R3 with 256
--											24 =>"0011100000000101",----------------------------LHI -Load R4 with 640
--											25 =>"0011101000000100",----------------------------LHI -Load R5 with 512
--											26 =>"0011110000000101",----------------------------LHI -Load R6 with 640
--											30 =>"0011111000000001",----------------------------LHI -Load R7 with 128
--											31 =>"1001000000001001",----------------------------JAL jump to 40 instruction 
--											32 =>"0011001000000000",-----------------------------LHI -Load R0 with 0
--											40 =>"0011000000000001",----------------------------LHI -Load R0 with 128
--											41 =>"1010001111000000",------------------------------JLR to 128
--											128 =>"0011111000000110",----------------------LHI -Load R7 with 768
--											129 =>"0011111000000000",----------------------LHI -Load R7 with 0
--											130 =>"1011000000001010",----------------------JRI to 138
--											138 =>"0011111000000110",----------------------LHI -Load R7 with 768
--											
                                 others=>(others => 'X'));

											
begin
process(read_ena,address,i_memory)
begin
instruction_out <= i_memory(to_integer(unsigned(address))); 
end process;
end Instruction_behave;

 